`timescale 1ns / 1ps


module dct_cordic_tb();
reg clk,rst;
reg [19:0]x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15;
wire [19:0]y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15;

dct_cordic dc1(clk,rst,x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,
y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15);

initial clk=1;
always #5 clk=~clk;

initial
begin
rst=1;
#100 rst=0;
x0=20'b0_0000010_0000_0000_0000;
x1=20'b0_0000010_0000_0000_0000;
x2=20'b0_0000011_0000_0000_0000;
x3=20'b0_0000100_0000_0000_0000;
x4=20'b0_0000101_0000_0000_0000;
x5=20'b0_0000110_0000_0000_0000;
x6=20'b0_0000111_0000_0000_0000;
x7=20'b0_0001000_0000_0000_0000;
x8=20'b0_0001001_0000_0000_0000;
x9=20'b0_0000001_1000_0000_0000;
x10=20'b0_0000010_1000_0000_0000;
x11=20'b0_0000011_1000_0000_0000;
x12=20'b0_0000100_1000_0000_0000;
x13=20'b0_0000101_1000_0000_0000;
x14=20'b0_0000110_1000_0000_0000;
x15=20'b0_0000111_1000_0000_0000;
end

endmodule
